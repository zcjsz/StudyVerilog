module ex_cnt(
    input   wire            sclk,  // 模拟晶振产生时钟
    input   wire            rst_n, // 模拟外部复位信号
    output  wire    [9:0]   cnt
);

    reg [9:0] cnt_r;

    always @(posedge sclk or negedge rst_n) begin
        if(rst_n == 1'b0)
            cnt_r <= 10'd0;
        else 
            cnt_r <= cnt_r + 1'b1;
    end

    assign cnt = cnt_r;


endmodule
